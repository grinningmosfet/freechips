magic
tech sky130A
magscale 1 2
timestamp 1681238406
<< metal1 >>
rect 12 149 74 330
rect 112 -202 170 62
rect 12 -461 74 -280
rect 208 -364 271 233
use sky130_fd_pr__nfet_01v8_EDB9KC *sky130_fd_pr__nfet_01v8_EDB9KC_0
timestamp 1681237416
transform 1 0 141 0 1 -322
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_M479BZ  sky130_fd_pr__pfet_01v8_M479BZ_0
timestamp 1681237537
transform 1 0 141 0 1 191
box -211 -261 211 261
<< labels >>
flabel metal1 12 149 74 330 0 FreeMono 160 90 0 0 VDD
port 1 nsew
flabel metal1 12 -461 74 -280 0 FreeMono 160 90 0 0 VSS
port 2 nsew
flabel metal1 112 -140 170 -34 0 FreeMono 160 0 0 0 I
port 3 nsew
flabel metal1 208 -140 271 -34 0 FreeMono 160 0 0 0 O
port 4 nsew
<< end >>
